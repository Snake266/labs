module ALU(
           input rst,
           input clk,
           input [31:0] A,
           input [31:0] B,
           input [2:0] F,

           output reg [31:0] Y
           );

endmodule // ALU
