module fifo(
            input  clk,
            input  rst,
            input  we,
            input  re,
            input  data_in,
            output data_out,
            output empty,
            output full
            );

endmodule // fifo
