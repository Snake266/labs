module main(
            input [9:0]  sw,
            input [1:0]  key,
            input        clk,
            output       ledr[9:0],
            output [6:0] hex0,
            output [6:0] hex1);


endmodule // main
