module transmitter(
                   input     clk,
                   input reg data,
                   input     start,
                   output    busy,
                   output    tx
                   );

   always @ (posedge clk or posedge clk) begin

   end

endmodule // transmitter
