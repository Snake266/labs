module transmitter(
                   input     clk,
                   input reg data,
                   input     start,
                   output    busy,
                   output    tx
                   );
   always @ (  ) begin

   end

endmodule // transmitter
