module DC2 (
            input [7:4] SW,
            output [4 : 0] OUT
            );
   assign OUT = SW;
endmodule // DC2
