module or32_bus(input a, b, output y);
   assign y = a | b;
endmodule // or32_bus
